LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;

ENTITY PIC IS
    GENERIC(ADDLOGIC :  STD_LOGIC_VECTOR(15 DOWNTO 0):=x"0C05";
            IR1ISR :    STD_LOGIC_VECTOR(15 DOWNTO 0):=x"0900";
            IR2ISR :    STD_LOGIC_VECTOR(15 DOWNTO 0):=x"0910";
            IR3ISR :    STD_LOGIC_VECTOR(15 DOWNTO 0):=x"0920"
            );
    PORT(
    IR1,IR2,IR3 :IN STD_LOGIC;
    ADDRBUS :IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    DATABUS :OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    INT :OUT STD_LOGIC
    );
END ENTITY;
ARCHITECTURE ARCH OF PIC IS
    TYPE MEMORY IS ARRAY(NATURAL RANGE<>) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL MEM:MEMORY(2 DOWNTO 0):=(IR3ISR,IR2ISR,IR1ISR);
BEGIN
    INT<='1' WHEN ((IR1 OR IR2 OR IR3)='1') ELSE '0';
    DATABUS<= MEM(0) WHEN (IR1='1' AND ADDRBUS=ADDLOGIC) ELSE MEM(1) WHEN (IR2='1' AND ADDRBUS=ADDLOGIC) ELSE MEM(2) WHEN (IR3='1' AND ADDRBUS=ADDLOGIC) ELSE (OTHERS=>'Z');
END ARCHITECTURE;
